interface and_if;
  
  logic input_a, input_b;
  logic output_y;
endinterface
