interface count_if #(parameter N);
 
  logic rst,clk;
  logic [N:0] counter;
  logic [N:0] counter_up; 
endinterface
