module top();

  
  and_intr inf();

 
  and_gate a1(inf);

  
  tb a2(inf);

endmodule 
